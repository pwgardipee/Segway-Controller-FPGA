module steer_en(clk,rst_n, lft_ld, rght_ld, en_steer, rider_off, ld_cell_diff);

  input clk;		    // 50MHz clock
  input rst_n;		    // Active low asynch reset
  input [11:0] lft_ld, rght_ld;    //Left and right load cells

  output reg en_steer;		// enables steering (goes to balance_cntrl)
  output reg rider_off;     // pulses high for one clock on transition back to initial state
  output [11:0] ld_cell_diff;	//Difference between left and right load cells


  wire diff_gt_eigth;	//Load cell difference is greater than 1/8 of total weight
  wire diff_gt_15_16;	//Load cell difference is greater than 15/16 of total weight
  wire sum_gt_min;		//True when total weight is greater than minimum required weight
  wire sum_lt_min;		//True when total weight is less than minimum required weight
  wire [11:0] intr_cell_diff;	//The difference between the left and right load cells
  wire [12:0] ld_sum;			//The sum of the left and right load cells
  wire tmr_full;				//High when timer is done counting

  reg [25:0] timer_cnt;			//Timer
  reg clr_tmr;				//Signal to clear timer

  localparam MIN_RIDER_WEIGHT = 12'h200;	//Min rider weight defined by project spec
  localparam HYSTERESIS = 6'h20;			//Used to avoid instability in case rider = min rider weight exactly
  parameter fast_sim = 0;					//Used to speed up simulation time

  //localparam IDLE = 2'b00;
  //localparam WAIT = 2'b01;
  //localparam STEER_EN = 2'b10;
  //reg [1:0] state, nxt_state;

  //Define states for state machines
  typedef enum reg [1:0] {IDLE, WAIT, STEER_EN} state_t;
  state_t state, nxt_state;

  //Sum of left and right load cells
  assign ld_sum = lft_ld + rght_ld;

  //Difference should be absolute value
  assign intr_cell_diff = (lft_ld > rght_ld) ? (lft_ld - rght_ld) : (rght_ld - lft_ld);

  //Assign output value
  assign ld_cell_diff = lft_ld - rght_ld;

  //Timer flip flop
  always_ff @(posedge clk, negedge rst_n)
    if(!rst_n)
	timer_cnt <= 26'h0000000;
    else if(clr_tmr)
	timer_cnt <= 26'h0000000;
    else
	timer_cnt <= timer_cnt + 1'b1;


	//Timer full based on 26 bit counter
	assign tmr_full = fast_sim ? &timer_cnt[14:0] : &timer_cnt;

	//diff_gt_eith = true when ld_cell_diff > 1/8*(left+right)
	assign diff_gt_eigth = (intr_cell_diff > ((ld_sum) >> 3));

	//diff_gt_15_16 = true when ld_cell_diff > 15/16(left + right)
	assign diff_gt_15_16 = (intr_cell_diff > ((ld_sum)-((ld_sum) >> 4)));

	//sum_gt_min = true when left+right > (min rider weight + hysteresis)
	assign sum_gt_min = ((ld_sum) > (MIN_RIDER_WEIGHT + HYSTERESIS));

	//sum_lt_min = true when  left+ right < (min rider weight - hysteresis)
	assign sum_lt_min = ((ld_sum) < (MIN_RIDER_WEIGHT - HYSTERESIS));

	//State Machine- Go to next state
	always_ff @(posedge clk, negedge rst_n)
	if(!rst_n)
		state <= IDLE;
	else
		state <= nxt_state;

always_comb begin

    en_steer = 1'b0;
    clr_tmr = 1'b0;
    nxt_state = IDLE;
    rider_off = 1'b0;
    case(state)
	IDLE:
			//Waiting for rider to put any weight on the segway
	    if(sum_gt_min) begin
		nxt_state = WAIT;
		clr_tmr = 1'b1;
	    end
	    else begin
		nxt_state = IDLE;
		rider_off = 1'b1;
	    end
	WAIT:
			//Waiting for rider to stabilize on the segway
	    if(!sum_gt_min) begin
				//Rider got off of segway
		nxt_state = IDLE;
		rider_off = 1'b1;
	    end
	    else if(diff_gt_eigth) begin
				//Rider is not stable yet
		nxt_state = WAIT;
		clr_tmr = 1'b1;
	    end
	    else if(tmr_full) begin
				//Rider is considered stable after 1.3 seconds
		nxt_state = STEER_EN;
		en_steer = 1'b1;
	    end
	    else
		nxt_state = WAIT;
	STEER_EN:
			//Steering is now enabled
	    if(sum_lt_min) begin
				//Rider is no longer on the segway
		nxt_state = IDLE;
		en_steer = 1'b0;
		rider_off = 1'b1;
	    end
	    else if(diff_gt_15_16) begin
				//Rider is no longer stable
		nxt_state = WAIT;
		clr_tmr = 1'b1;
		en_steer = 1'b0;
	    end
	    else if(!diff_gt_15_16) begin
				//Rider is still stable
		en_steer = 1'b1;
		nxt_state = STEER_EN;
	    end
	    else
		nxt_state = STEER_EN;
    endcase

end

endmodule
